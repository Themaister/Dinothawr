BSV1                                                                                                                        